VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ms00f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN ck DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END ck
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.05 0.500 1.15 1.500 ;
    END
  END d
END ms00f80

MACRO oa22f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END oa22f80

MACRO oa22f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END oa22f40

MACRO oa22f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END oa22f20

MACRO oa22f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END oa22f10

MACRO oa22f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END oa22f08

MACRO oa22f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END oa22f06

MACRO oa22f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END oa22f04

MACRO oa22f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END oa22f03

MACRO oa22f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END oa22f02

MACRO oa22f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN d 
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END d
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN o 
    TAPERRULE EM_NDR ;
    DIRECTION OUTPUT ;
    PORT
    LAYER metal2 ;  
      RECT 1.25 0.500 1.35 1.050 ;
      RECT 1.35 0.950 1.55 1.050 ;
    END
  END o
END oa22f01

MACRO oa22m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END oa22m80

MACRO oa22m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END oa22m40

MACRO oa22m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END oa22m20

MACRO oa22m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END oa22m10

MACRO oa22m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END oa22m08

MACRO oa22m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END oa22m06

MACRO oa22m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END oa22m04

MACRO oa22m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END oa22m03

MACRO oa22m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END oa22m02

MACRO oa22m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END oa22m01

MACRO oa22s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END oa22s80

MACRO oa22s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END oa22s40

MACRO oa22s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END oa22s20

MACRO oa22s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END oa22s10

MACRO oa22s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END oa22s08

MACRO oa22s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END oa22s06

MACRO oa22s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END oa22s04

MACRO oa22s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END oa22s03

MACRO oa22s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END oa22s02

MACRO oa22s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END oa22s01

MACRO oa12f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END oa12f80

MACRO oa12f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END oa12f40

MACRO oa12f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END oa12f20

MACRO oa12f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END oa12f10

MACRO oa12f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END oa12f08

MACRO oa12f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END oa12f06

MACRO oa12f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END oa12f04

MACRO oa12f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END oa12f03

MACRO oa12f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END oa12f02

MACRO oa12f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END oa12f01

MACRO oa12m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END oa12m80

MACRO oa12m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END oa12m40

MACRO oa12m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END oa12m20

MACRO oa12m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END oa12m10

MACRO oa12m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END oa12m08

MACRO oa12m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END oa12m06

MACRO oa12m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END oa12m04

MACRO oa12m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END oa12m03

MACRO oa12m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END oa12m02

MACRO oa12m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END oa12m01

MACRO oa12s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END oa12s80

MACRO oa12s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END oa12s40

MACRO oa12s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END oa12s20

MACRO oa12s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END oa12s10

MACRO oa12s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END oa12s08

MACRO oa12s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END oa12s06

MACRO oa12s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END oa12s04

MACRO oa12s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END oa12s03

MACRO oa12s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END oa12s02

MACRO oa12s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END oa12s01

MACRO ao22f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END ao22f80

MACRO ao22f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END ao22f40

MACRO ao22f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END ao22f20

MACRO ao22f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END ao22f10

MACRO ao22f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END ao22f08

MACRO ao22f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END ao22f06

MACRO ao22f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END ao22f04

MACRO ao22f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END ao22f03

MACRO ao22f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END ao22f02

MACRO ao22f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END ao22f01

MACRO ao22m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END ao22m80

MACRO ao22m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END ao22m40

MACRO ao22m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END ao22m20

MACRO ao22m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END ao22m10

MACRO ao22m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END ao22m08

MACRO ao22m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END ao22m06

MACRO ao22m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END ao22m04

MACRO ao22m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END ao22m03

MACRO ao22m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END ao22m02

MACRO ao22m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END ao22m01

MACRO ao22s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 204.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 122.8 0.500 122.9 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 163.9 0.500 164 1.500 ;
    END
  END d
END ao22s80

MACRO ao22s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 61.45 0.500 61.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 81.85 0.500 81.95 1.500 ;
    END
  END d
END ao22s40

MACRO ao22s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 30.65 0.500 30.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 40.85 0.500 40.95 1.500 ;
    END
  END d
END ao22s20

MACRO ao22s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 15.25 0.500 15.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 20.45 0.500 20.55 1.500 ;
    END
  END d
END ao22s10

MACRO ao22s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 10.25 0.500 10.35 1.500 ;
    END
  END d
END ao22s08

MACRO ao22s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.65 0.500 5.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.65 0.500 7.75 1.500 ;
    END
  END d
END ao22s06

MACRO ao22s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END ao22s04

MACRO ao22s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.85 0.500 2.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END d
END ao22s03

MACRO ao22s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END ao22s02

MACRO ao22s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 1 ;
    EDGETYPE RIGHT 2 ;
  " ;

  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END ao22s01

MACRO ao12f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END ao12f80

MACRO ao12f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END ao12f40

MACRO ao12f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END ao12f20

MACRO ao12f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END ao12f10

MACRO ao12f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END ao12f08

MACRO ao12f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END ao12f06

MACRO ao12f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END ao12f04

MACRO ao12f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END ao12f03

MACRO ao12f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END ao12f02

MACRO ao12f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END ao12f01

MACRO ao12m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END ao12m80

MACRO ao12m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END ao12m40

MACRO ao12m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END ao12m20

MACRO ao12m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END ao12m10

MACRO ao12m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END ao12m08

MACRO ao12m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END ao12m06

MACRO ao12m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END ao12m04

MACRO ao12m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END ao12m03

MACRO ao12m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END ao12m02

MACRO ao12m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END ao12m01

MACRO ao12s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 153.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 115.2 0.500 115.3 1.500 ;
    END
  END c
END ao12s80

MACRO ao12s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 57.65 0.500 57.75 1.500 ;
    END
  END c
END ao12s40

MACRO ao12s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 28.85 0.500 28.95 1.500 ;
    END
  END c
END ao12s20

MACRO ao12s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 14.45 0.500 14.55 1.500 ;
    END
  END c
END ao12s10

MACRO ao12s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 7.25 0.500 7.35 1.500 ;
    END
  END c
END ao12s08

MACRO ao12s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 7.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.45 0.500 5.55 1.500 ;
    END
  END c
END ao12s06

MACRO ao12s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END ao12s04

MACRO ao12s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END ao12s03

MACRO ao12s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END ao12s02

MACRO ao12s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END ao12s01

MACRO no04f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END no04f80

MACRO no04f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END no04f40

MACRO no04f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END no04f20

MACRO no04f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END no04f10

MACRO no04f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END no04f08

MACRO no04f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END no04f06

MACRO no04f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END no04f04

MACRO no04f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END no04f03

MACRO no04f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END no04f02

MACRO no04f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END no04f01

MACRO no04m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END no04m80

MACRO no04m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END no04m40

MACRO no04m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END no04m20

MACRO no04m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END no04m10

MACRO no04m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END no04m08

MACRO no04m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END no04m06

MACRO no04m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END no04m04

MACRO no04m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END no04m03

MACRO no04m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END no04m02

MACRO no04m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END no04m01

MACRO no04s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END no04s80

MACRO no04s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END no04s40

MACRO no04s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END no04s20

MACRO no04s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END no04s10

MACRO no04s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END no04s08

MACRO no04s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END no04s06

MACRO no04s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END no04s04

MACRO no04s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END no04s03

MACRO no04s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END no04s02

MACRO no04s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END no04s01

MACRO no03f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END no03f80

MACRO no03f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END no03f40

MACRO no03f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END no03f20

MACRO no03f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END no03f10

MACRO no03f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END no03f08

MACRO no03f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END no03f06

MACRO no03f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END no03f04

MACRO no03f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END no03f03

MACRO no03f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END no03f02

MACRO no03f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END no03f01

MACRO no03m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END no03m80

MACRO no03m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END no03m40

MACRO no03m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END no03m20

MACRO no03m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END no03m10

MACRO no03m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END no03m08

MACRO no03m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END no03m06

MACRO no03m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END no03m04

MACRO no03m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END no03m03

MACRO no03m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END no03m02

MACRO no03m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END no03m01

MACRO no03s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END no03s80

MACRO no03s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END no03s40

MACRO no03s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END no03s20

MACRO no03s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END no03s10

MACRO no03s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END no03s08

MACRO no03s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END no03s06

MACRO no03s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END no03s04

MACRO no03s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END no03s03

MACRO no03s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END no03s02

MACRO no03s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END no03s01

MACRO no02f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END no02f80

MACRO no02f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END no02f40

MACRO no02f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END no02f20

MACRO no02f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END no02f10

MACRO no02f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END no02f08

MACRO no02f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END no02f06

MACRO no02f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END no02f04

MACRO no02f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END no02f03

MACRO no02f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END no02f02

MACRO no02f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END no02f01

MACRO no02m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END no02m80

MACRO no02m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END no02m40

MACRO no02m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END no02m20

MACRO no02m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END no02m10

MACRO no02m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END no02m08

MACRO no02m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END no02m06

MACRO no02m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END no02m04

MACRO no02m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END no02m03

MACRO no02m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END no02m02

MACRO no02m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END no02m01

MACRO no02s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END no02s80

MACRO no02s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END no02s40

MACRO no02s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END no02s20

MACRO no02s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END no02s10

MACRO no02s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END no02s08

MACRO no02s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END no02s06

MACRO no02s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END no02s04

MACRO no02s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END no02s03

MACRO no02s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END no02s02

MACRO no02s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END no02s01

MACRO na04f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END na04f80

MACRO na04f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END na04f40

MACRO na04f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END na04f20

MACRO na04f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END na04f10

MACRO na04f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END na04f08

MACRO na04f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END na04f06

MACRO na04f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END na04f04

MACRO na04f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END na04f03

MACRO na04f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END na04f02

MACRO na04f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END na04f01

MACRO na04m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END na04m80

MACRO na04m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END na04m40

MACRO na04m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END na04m20

MACRO na04m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END na04m10

MACRO na04m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END na04m08

MACRO na04m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END na04m06

MACRO na04m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END na04m04

MACRO na04m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END na04m03

MACRO na04m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END na04m02

MACRO na04m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END na04m01

MACRO na04s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 128.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 102.5 0.500 102.6 1.500 ;
    END
  END d
END na04s80

MACRO na04s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 64.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.45 0.500 38.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END d
END na04s40

MACRO na04s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 32.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END d
END na04s20

MACRO na04s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 16.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.65 0.500 9.75 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END d
END na04s10

MACRO na04s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 8.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END d
END na04s08

MACRO na04s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.85 0.500 3.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 5.05 0.500 5.15 1.500 ;
    END
  END d
END na04s06

MACRO na04s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END d
END na04s04

MACRO na04s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END d
END na04s03

MACRO na04s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.45 0.500 1.55 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END d
END na04s02

MACRO na04s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
  PIN d DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END d
END na04s01

MACRO na03f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END na03f80

MACRO na03f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END na03f40

MACRO na03f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END na03f20

MACRO na03f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END na03f10

MACRO na03f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END na03f08

MACRO na03f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END na03f06

MACRO na03f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END na03f04

MACRO na03f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END na03f03

MACRO na03f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END na03f02

MACRO na03f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END na03f01

MACRO na03m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END na03m80

MACRO na03m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END na03m40

MACRO na03m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END na03m20

MACRO na03m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END na03m10

MACRO na03m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END na03m08

MACRO na03m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END na03m06

MACRO na03m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END na03m04

MACRO na03m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END na03m03

MACRO na03m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END na03m02

MACRO na03m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END na03m01

MACRO na03s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 102.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 76.85 0.500 76.95 1.500 ;
    END
  END c
END na03s80

MACRO na03s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.85 0.500 25.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 38.65 0.500 38.75 1.500 ;
    END
  END c
END na03s40

MACRO na03s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 19.25 0.500 19.35 1.500 ;
    END
  END c
END na03s20

MACRO na03s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 13.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.65 0.500 6.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 9.85 0.500 9.95 1.500 ;
    END
  END c
END na03s10

MACRO na03s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 4.85 0.500 4.95 1.500 ;
    END
  END c
END na03s08

MACRO na03s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.65 0.500 3.75 1.500 ;
    END
  END c
END na03s06

MACRO na03s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.65 0.500 2.75 1.500 ;
    END
  END c
END na03s04

MACRO na03s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.85 0.500 1.95 1.500 ;
    END
  END c
END na03s03

MACRO na03s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END c
END na03s02

MACRO na03s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END b
  PIN c DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END c
END na03s01

MACRO na02f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END na02f80

MACRO na02f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END na02f40

MACRO na02f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END na02f20

MACRO na02f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END na02f10

MACRO na02f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END na02f08

MACRO na02f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END na02f06

MACRO na02f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END na02f04

MACRO na02f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END na02f03

MACRO na02f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END na02f02

MACRO na02f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END na02f01

MACRO na02m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END na02m80

MACRO na02m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END na02m40

MACRO na02m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END na02m20

MACRO na02m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END na02m10

MACRO na02m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END na02m08

MACRO na02m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END na02m06

MACRO na02m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END na02m04

MACRO na02m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END na02m03

MACRO na02m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END na02m02

MACRO na02m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END na02m01

MACRO na02s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 76.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 51.25 0.500 51.35 1.500 ;
    END
  END b
END na02s80

MACRO na02s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 38.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END b
END na02s40

MACRO na02s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 19.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END b
END na02s20

MACRO na02s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 9.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END b
END na02s10

MACRO na02s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 4.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END b
END na02s08

MACRO na02s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 2.45 0.500 2.55 1.500 ;
    END
  END b
END na02s06

MACRO na02s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END b
END na02s04

MACRO na02s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.0 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END b
END na02s03

MACRO na02s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END b
END na02s02

MACRO na02s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
  PIN b DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END b
END na02s01

MACRO in01f80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
END in01f80

MACRO in01f40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
END in01f40

MACRO in01f20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
END in01f20

MACRO in01f10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
END in01f10

MACRO in01f08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
END in01f08

MACRO in01f06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
END in01f06

MACRO in01f04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
END in01f04

MACRO in01f03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
END in01f03

MACRO in01f02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
END in01f02

MACRO in01f01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
#       LAYER metal2 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
END in01f01

MACRO in01m80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
END in01m80

MACRO in01m40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
END in01m40

MACRO in01m20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
END in01m20

MACRO in01m10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
END in01m10

MACRO in01m08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
END in01m08

MACRO in01m06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
END in01m06

MACRO in01m04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
END in01m04

MACRO in01m03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
END in01m03

MACRO in01m02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
END in01m02

MACRO in01m01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
END in01m01

MACRO in01s80
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 51.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 25.65 0.500 25.75 1.500 ;
    END
  END a
END in01s80

MACRO in01s40
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 25.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 12.85 0.500 12.95 1.500 ;
    END
  END a
END in01s40

MACRO in01s20
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 12.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 6.45 0.500 6.55 1.500 ;
    END
  END a
END in01s20

MACRO in01s10
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END a
END in01s10

MACRO in01s08
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 3.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.65 0.500 1.75 1.500 ;
    END
  END a
END in01s08

MACRO in01s06
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 2.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 1.25 0.500 1.35 1.500 ;
    END
  END a
END in01s06

MACRO in01s04
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END a
END in01s04

MACRO in01s03
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.65 0.500 0.75 1.500 ;
    END
  END a
END in01s03

MACRO in01s02
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END a
END in01s02

MACRO in01s01
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.4 BY 2.0 ;
  SYMMETRY X Y R90 ;

  SITE  core ;
  PIN o DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END o
  PIN a DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.25 0.500 0.35 1.500 ;
    END
  END a
END in01s01

MACRO b
     SIZE 300.000 BY 200.0 ;
     ORIGIN 0 0 ;
     SYMMETRY X Y ;
     SITE core ;
     CLASS BLOCK ;  
     PIN i1 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 0.00 0.000 1.00 1.00 ;
      END
     END i1
     PIN i2 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 5.00 0.000 6.0 1.00 ;
      END
     END i2
     PIN i3 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 10.0 0.000 11.00 1.000 ;
      END
     END i3
     PIN i4 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 15.00 0.00 16.00 1.000 ;
      END
     END i4
     PIN i5 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 20.0 0.00 21.0 1.00 ;
      END
     END i5
     PIN i6 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 30.0 0.00 31.0 1.00 ;
      END
     END i6
     PIN i7 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 35.0 0.00 36.0 1.00 ;
      END
     END i7
     PIN i8 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 40.0 0.00 41.0 1.00 ;
      END
     END i8
     PIN i9 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 45.0 0.00 46.0 1.00 ;
      END
     END i9
     PIN i10 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 50.0 0.00 51.0 1.00 ;
      END
     END i10
     PIN i11 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 55.0 0.00 56.0 1.00 ;
      END
     END i11
     PIN i12 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 60.0 0.00 61.0 1.00 ;
      END
     END i12
     PIN i13 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 65.0 0.00 66.0 1.00 ;
      END
     END i13
     PIN i14 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 70.0 0.00 71.0 1.00 ;
      END
     END i14
     PIN i15 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 75.0 0.00 76.0 1.00 ;
      END
     END i15
     PIN i16 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 80.0 0.00 81.0 1.00 ;
      END
     END i16
     PIN i17 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 85.0 0.00 86.0 1.00 ;
      END
     END i17
     PIN i18 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 90.0 0.00 91.0 1.00 ;
      END
     END i18
     PIN i19 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 95.0 0.00 96.0 1.00 ;
      END
     END i19
     PIN i20 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 100.0 0.00 101.0 1.00 ;
      END
     END i20
     OBS 
          LAYER metal1 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal2 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal3 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal4 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
END b

MACRO c
     SIZE 300.000 BY 200.0 ;
     ORIGIN 0 0 ;
     SYMMETRY X Y ;
     SITE core ;
     CLASS BLOCK ;  
     PIN i1 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 0.00 0.000 1.00 1.00 ;
      END
     END i1
     PIN i2 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 5.00 0.000 6.0 1.00 ;
      END
     END i2
     PIN i3 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 10.0 0.000 11.00 1.000 ;
      END
     END i3
     PIN i4 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 15.00 0.00 16.00 1.000 ;
      END
     END i4
     PIN i5 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 20.0 0.00 21.0 1.00 ;
      END
     END i5
     PIN i6 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 25.0 0.00 26.0 1.00 ;
      END
     END i6
     PIN i7 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 35.0 0.00 36.0 1.00 ;
      END
     END i7
     PIN i8 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 40.0 0.00 41.0 1.00 ;
      END
     END i8
     PIN i9 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 45.0 0.00 46.0 1.00 ;
      END
     END i9
     PIN i10 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 50.0 0.00 51.0 1.00 ;
      END
     END i10
     PIN i11 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 55.0 0.00 56.0 1.00 ;
      END
     END i11
     PIN i12 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 60.0 0.00 61.0 1.00 ;
      END
     END i12
     PIN i13 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 65.0 0.00 66.0 1.00 ;
      END
     END i13
     PIN i14 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 70.0 0.00 71.0 1.00 ;
      END
     END i14
     PIN i15 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 75.0 0.00 76.0 1.00 ;
      END
     END i15
     PIN i16 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 80.0 0.00 81.0 1.00 ;
      END
     END i16
     PIN i17 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 85.0 0.00 86.0 1.00 ;
      END
     END i17
     PIN i18 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 90.0 0.00 91.0 1.00 ;
      END
     END i18
     PIN i19 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 95.0 0.00 96.0 1.00 ;
      END
     END i19
     PIN i20 DIRECTION INPUT ;
      PORT
        LAYER metal1 ;
        RECT 100.0 0.00 101.0 1.00 ;
      END
     END i20
     OBS 
          LAYER metal1 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal2 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal3 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
     OBS 
          LAYER metal4 ;
               RECT 0.000 0.000 300.000 200.000 ;
     END
END c

END LIBRARY

END LIBRARY
